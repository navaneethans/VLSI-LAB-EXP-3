module ha(a,b,sum,carry);
input a,b;
output sum,carry;

endmodule

module multi_2(a,b,p,carry);
input [1:0]a,b;
output [2:0]p;
output carry;

endmodule
