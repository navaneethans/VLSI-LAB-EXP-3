module ha(a,b,sum,carry);
input a,b;
output sum,carry;


endmodule

module fa_ha(a,b,c,sum,carry);
input a,b,c;
output sum,carry;


endmodule

module multi_4(a,b,p,carry);
input[3:0]a,b;
output [6:0]p;
output carry;
wire [17:1]w;




endmodule
